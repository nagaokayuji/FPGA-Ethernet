/*
control to byte_data

*/

module send_control(

)